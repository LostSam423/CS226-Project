library ieee;
use ieee.std_logic_1164.all;

entity DFlipFlop is
	port (clk, rst, d: in std_logic; s: out std_logic);
end entity;

architecture behave of DFlipFlop is
begin
	process (clk)
	begin
		if (rising_edge(clk)) then
			if (rst = '1' ) then
				s <= '0';
			else
				s <= d;
			end if;
		end if;
	end process;
end architecture;